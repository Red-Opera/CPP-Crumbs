0 0 0 0 0 0                                                                                          0 0 0 0 0 0                                                                                          0 0 0 0 0 0                                                                                          0 0 0 0 0 00000000000000000000000000000000000000000000000000000000000000000000000000000000000 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 2 2 0 0 0 0 